module ESM_core (
    input [31:0] Instr_in,
    output reg [3:0]Buffer_index 
);
    
endmodule